module memory(clk,rst,wt_rd,addr,wdata,rdata,valid,ready);
parameter WIDTH=16;
parameter DEPTH=64;
parameter ADDR_WIDTH=$clog2(DEPTH);

input clk,rst;
input wt_rd;
input [ADDR_WIDTH-1:0]addr;
input [WIDTH-1:0]wdata;
output reg [WIDTH-1:0]rdata;
input valid;
output reg ready;
integer i;

reg [WIDTH-1:0] mem [DEPTH-1:0];

always@(posedge clk) begin
	if(rst) begin
		rdata=0;
		ready=0;
		for(i=0;i<DEPTH;i=i+1) begin
			mem[i]=0;
		end
	end
	else begin
		if(valid) begin
			ready=1;
			if(wt_rd) begin
				mem[addr]=wdata;
			end
			else begin
				rdata=mem[addr];
			end
		end
		else begin
			ready=0;
		end
	end
end

endmodule
