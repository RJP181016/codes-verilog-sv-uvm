module top;
reg clk,rst;
mem_common mem_common_i=new();

//DUT instance
memory #(.WIDTH(`WIDTH),.DEPTH(`DEPTH),.ADDR_WIDTH(`ADDR_WIDTH)) dut (.clk(pif.clk),
			.rst(pif.rst),
			.wt_rd(pif.wt_rd),
			.addr(pif.addr),
			.wdata(pif.wdata),
			.rdata(pif.rdata),
			.valid(pif.valid),
			.ready(pif.ready)
			);
//clk gen
initial begin
	clk=0;
	forever #5 clk = ~clk;
end

mem_env env;
//reset
initial begin
	rst=0;
	#5;
	rst=1;
	reset_mem();
	#20;
	rst=0;

	env=new();
	env.run();
end

//interface instance
mem_intf pif(clk,rst);

initial begin
mem_common::vif=pif;
end




task reset_mem();
	pif.addr=0;
	pif.wdata=0;
	pif.valid=0;
	pif.wt_rd=0;
endtask

initial begin
	$value$plusargs("testname=%s",mem_common::testname);
	wait(mem_common::count*2*mem_common::num_agents==mem_common::total_tx_driven);
	#20;
	if(mem_common::num_mismatches!=0 || mem_common::num_matches!=mem_common::num_agents*mem_common::count) begin
		$display("#### TEST FAILED ####");
		$display("## num_matches=%0d ##",mem_common::num_matches);
		$display("## num_mismatches=%0d ##",mem_common::num_mismatches);
	end
	else $display("#### TEST PASSED ####");
	$display("addr_width",`ADDR_WIDTH);
	$finish;
end

endmodule
