`include "dma_axi64.v"
`include "dma_axi64_apb_mux.v"
`include "dma_axi64_ch_reg_params.v"
`include "dma_axi64_core0.v"
`include "dma_axi64_core0_arbiter.v"
`include "dma_axi64_core0_axim_cmd.v"
`include "dma_axi64_core0_axim_rd.v"
`include "dma_axi64_core0_axim_rdata.v"
`include "dma_axi64_core0_axim_resp.v"
`include "dma_axi64_core0_axim_timeout.v"
`include "dma_axi64_core0_axim_wdata.v"
`include "dma_axi64_core0_axim_wr.v"
`include "dma_axi64_core0_ch.v"
`include "dma_axi64_core0_ch_calc.v"
`include "dma_axi64_core0_ch_calc_addr.v"
`include "dma_axi64_core0_ch_calc_joint.v"
`include "dma_axi64_core0_ch_calc_size.v"
//`include "dma_axi64_core0_ch_empty.v"
`include "dma_axi64_core0_ch_fifo.v"
`include "dma_axi64_core0_ch_fifo_ctrl.v"
`include "dma_axi64_core0_ch_fifo_ptr.v"
`include "dma_axi64_core0_ch_offsets.v"
`include "dma_axi64_core0_ch_outs.v"
`include "dma_axi64_core0_ch_periph_mux.v"
`include "dma_axi64_core0_ch_rd_slicer.v"
`include "dma_axi64_core0_ch_reg.v"
`include "dma_axi64_core0_ch_reg_size.v"
`include "dma_axi64_core0_ch_remain.v"
`include "dma_axi64_core0_ch_wr_slicer.v"
`include "dma_axi64_core0_channels.v"
`include "dma_axi64_core0_channels_apb_mux.v"
`include "dma_axi64_core0_channels_mux.v"
`include "dma_axi64_core0_ctrl.v"
`include "dma_axi64_core0_top.v"
`include "dma_axi64_core0_wdt.v"
`include "dma_axi64_defines.v"
`include "dma_axi64_dual_core.v"
`include "dma_axi64_reg.v"
`include "dma_axi64_reg_core0.v"
`include "dma_axi64_reg_params.v"
`include "prgen_delay.v"
`include "prgen_demux8.v"
`include "prgen_fifo.v"
`include "prgen_joint_stall.v"
`include "prgen_min2.v"
`include "prgen_min3.v"
`include "prgen_mux8.v"
`include "prgen_or8.v"
`include "prgen_rawstat.v"
`include "prgen_scatter8_1.v"
`include "prgen_stall.v"
`include "prgen_swap_32.v"
`include "prgen_swap_64.v"

