class eth_common;
//static mailbox gen2bfm=new();
static int pkt_count=10;
endclass
