register write read test
	STATIC_REG3 is not implemented in design
