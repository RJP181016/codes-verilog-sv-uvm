`include "uvm_macros.svh"
import uvm_pkg::*;

`include "packet.sv"
`include "test.sv"

program test;
  
  initial run_test();
  
endprogram
