`include "uvm_macros.svh"
import uvm_pkg::*;

`include "write_tx.sv"
`include "read_tx.sv"
`include "write_seq_lib.sv"
`include "read_seq_lib.sv"
`include "write_drv.sv"
`include "read_drv.sv"
`include "write_sqr.sv"
`include "read_sqr.sv"
`include "write_mon.sv"
`include "read_mon.sv"
`include "write_cov.sv"
`include "read_cov.sv"
`include "fifo_sbd.sv"
`include "write_agent.sv"
`include "read_agent.sv"
`include "fifo_env.sv"
`include "test_lib.sv"
