class apb_cov extends uvm_subscriber#(apb_tx);
`uvm_component_utils(apb_cov)
apb_tx tx;

covergroup apb_cg;
	ADDR_CP: coverpoint tx.addr {
		bins CH0_CMD_REG0 = {`CH0_CMD_REG0_ADDR};
        bins CH0_CMD_REG1 = {`CH0_CMD_REG1_ADDR};
        bins CH0_CMD_REG2 = {`CH0_CMD_REG2_ADDR};
        bins CH0_CMD_REG3 = {`CH0_CMD_REG3_ADDR};
        bins CH0_STATIC_REG0 = {`CH0_STATIC_REG0_ADDR};
        bins CH0_STATIC_REG1 = {`CH0_STATIC_REG1_ADDR};
        bins CH0_STATIC_REG2 = {`CH0_STATIC_REG2_ADDR};
        bins CH0_STATIC_REG3 = {`CH0_STATIC_REG3_ADDR};
        bins CH0_STATIC_REG4 = {`CH0_STATIC_REG4_ADDR};
        bins CH0_RESTRICT_REG = {`CH0_RESTRICT_REG_ADDR};
        bins CH0_READ_OFFSET_REG = {`CH0_READ_OFFSET_REG_ADDR};
        bins CH0_WRITE_OFFSET_REG = {`CH0_WRITE_OFFSET_REG_ADDR};
        bins CH0_FIFO_FULLNESS_REG = {`CH0_FIFO_FULLNESS_REG_ADDR};
        bins CH0_CMD_OUTS_REG = {`CH0_CMD_OUTS_REG_ADDR};
        bins CH0_CH_ENABLE_REG = {`CH0_CH_ENABLE_REG_ADDR};
        bins CH0_CH_START_REG = {`CH0_CH_START_REG_ADDR};
        bins CH0_CH_ACTIVE_REG = {`CH0_CH_ACTIVE_REG_ADDR};
        bins CH0_COUNT_REG = {`CH0_COUNT_REG_ADDR};
        bins CH0_INT_RAWSTAT_REG = {`CH0_INT_RAWSTAT_REG_ADDR};
        bins CH0_INT_CLEAR_REG = {`CH0_INT_CLEAR_REG_ADDR};
        bins CH0_INT_ENABLE_REG = {`CH0_INT_ENABLE_REG_ADDR};
        bins CH0_INT_STATUS_REG = {`CH0_INT_STATUS_REG_ADDR};
        bins CH1_CMD_REG0 = {`CH1_CMD_REG0_ADDR};
        bins CH1_CMD_REG1 = {`CH1_CMD_REG1_ADDR};
        bins CH1_CMD_REG2 = {`CH1_CMD_REG2_ADDR};
        bins CH1_CMD_REG3 = {`CH1_CMD_REG3_ADDR};
        bins CH1_STATIC_REG0 = {`CH1_STATIC_REG0_ADDR};
        bins CH1_STATIC_REG1 = {`CH1_STATIC_REG1_ADDR};
        bins CH1_STATIC_REG2 = {`CH1_STATIC_REG2_ADDR};
        bins CH1_STATIC_REG3 = {`CH1_STATIC_REG3_ADDR};
        bins CH1_STATIC_REG4 = {`CH1_STATIC_REG4_ADDR};
        bins CH1_RESTRICT_REG = {`CH1_RESTRICT_REG_ADDR};
        bins CH1_READ_OFFSET_REG = {`CH1_READ_OFFSET_REG_ADDR};
        bins CH1_WRITE_OFFSET_REG = {`CH1_WRITE_OFFSET_REG_ADDR};
        bins CH1_FIFO_FULLNESS_REG = {`CH1_FIFO_FULLNESS_REG_ADDR};
        bins CH1_CMD_OUTS_REG = {`CH1_CMD_OUTS_REG_ADDR};
        bins CH1_CH_ENABLE_REG = {`CH1_CH_ENABLE_REG_ADDR};
        bins CH1_CH_START_REG = {`CH1_CH_START_REG_ADDR};
        bins CH1_CH_ACTIVE_REG = {`CH1_CH_ACTIVE_REG_ADDR};
        bins CH1_COUNT_REG = {`CH1_COUNT_REG_ADDR};
        bins CH1_INT_RAWSTAT_REG = {`CH1_INT_RAWSTAT_REG_ADDR};
        bins CH1_INT_CLEAR_REG = {`CH1_INT_CLEAR_REG_ADDR};
        bins CH1_INT_ENABLE_REG = {`CH1_INT_ENABLE_REG_ADDR};
        bins CH1_INT_STATUS_REG = {`CH1_INT_STATUS_REG_ADDR};
        bins CH2_CMD_REG0 = {`CH2_CMD_REG0_ADDR};
        bins CH2_CMD_REG1 = {`CH2_CMD_REG1_ADDR};
        bins CH2_CMD_REG2 = {`CH2_CMD_REG2_ADDR};
        bins CH2_CMD_REG3 = {`CH2_CMD_REG3_ADDR};
        bins CH2_STATIC_REG0 = {`CH2_STATIC_REG0_ADDR};
        bins CH2_STATIC_REG1 = {`CH2_STATIC_REG1_ADDR};
        bins CH2_STATIC_REG2 = {`CH2_STATIC_REG2_ADDR};
        bins CH2_STATIC_REG3 = {`CH2_STATIC_REG3_ADDR};
        bins CH2_STATIC_REG4 = {`CH2_STATIC_REG4_ADDR};
        bins CH2_RESTRICT_REG = {`CH2_RESTRICT_REG_ADDR};
        bins CH2_READ_OFFSET_REG = {`CH2_READ_OFFSET_REG_ADDR};
        bins CH2_WRITE_OFFSET_REG = {`CH2_WRITE_OFFSET_REG_ADDR};
        bins CH2_FIFO_FULLNESS_REG = {`CH2_FIFO_FULLNESS_REG_ADDR};
        bins CH2_CMD_OUTS_REG = {`CH2_CMD_OUTS_REG_ADDR};
        bins CH2_CH_ENABLE_REG = {`CH2_CH_ENABLE_REG_ADDR};
        bins CH2_CH_START_REG = {`CH2_CH_START_REG_ADDR};
        bins CH2_CH_ACTIVE_REG = {`CH2_CH_ACTIVE_REG_ADDR};
        bins CH2_COUNT_REG = {`CH2_COUNT_REG_ADDR};
        bins CH2_INT_RAWSTAT_REG = {`CH2_INT_RAWSTAT_REG_ADDR};
        bins CH2_INT_CLEAR_REG = {`CH2_INT_CLEAR_REG_ADDR};
        bins CH2_INT_ENABLE_REG = {`CH2_INT_ENABLE_REG_ADDR};
        bins CH2_INT_STATUS_REG = {`CH2_INT_STATUS_REG_ADDR};
        bins CH3_CMD_REG0 = {`CH3_CMD_REG0_ADDR};
        bins CH3_CMD_REG1 = {`CH3_CMD_REG1_ADDR};
        bins CH3_CMD_REG2 = {`CH3_CMD_REG2_ADDR};
        bins CH3_CMD_REG3 = {`CH3_CMD_REG3_ADDR};
        bins CH3_STATIC_REG0 = {`CH3_STATIC_REG0_ADDR};
        bins CH3_STATIC_REG1 = {`CH3_STATIC_REG1_ADDR};
        bins CH3_STATIC_REG2 = {`CH3_STATIC_REG2_ADDR};
        bins CH3_STATIC_REG3 = {`CH3_STATIC_REG3_ADDR};
        bins CH3_STATIC_REG4 = {`CH3_STATIC_REG4_ADDR};
        bins CH3_RESTRICT_REG = {`CH3_RESTRICT_REG_ADDR};
        bins CH3_READ_OFFSET_REG = {`CH3_READ_OFFSET_REG_ADDR};
        bins CH3_WRITE_OFFSET_REG = {`CH3_WRITE_OFFSET_REG_ADDR};
        bins CH3_FIFO_FULLNESS_REG = {`CH3_FIFO_FULLNESS_REG_ADDR};
        bins CH3_CMD_OUTS_REG = {`CH3_CMD_OUTS_REG_ADDR};
        bins CH3_CH_ENABLE_REG = {`CH3_CH_ENABLE_REG_ADDR};
        bins CH3_CH_START_REG = {`CH3_CH_START_REG_ADDR};
        bins CH3_CH_ACTIVE_REG = {`CH3_CH_ACTIVE_REG_ADDR};
        bins CH3_COUNT_REG = {`CH3_COUNT_REG_ADDR};
        bins CH3_INT_RAWSTAT_REG = {`CH3_INT_RAWSTAT_REG_ADDR};
        bins CH3_INT_CLEAR_REG = {`CH3_INT_CLEAR_REG_ADDR};
        bins CH3_INT_ENABLE_REG = {`CH3_INT_ENABLE_REG_ADDR};
        bins CH3_INT_STATUS_REG = {`CH3_INT_STATUS_REG_ADDR};
        bins CH4_CMD_REG0 = {`CH4_CMD_REG0_ADDR};
        bins CH4_CMD_REG1 = {`CH4_CMD_REG1_ADDR};
        bins CH4_CMD_REG2 = {`CH4_CMD_REG2_ADDR};
        bins CH4_CMD_REG3 = {`CH4_CMD_REG3_ADDR};
        bins CH4_STATIC_REG0 = {`CH4_STATIC_REG0_ADDR};
        bins CH4_STATIC_REG1 = {`CH4_STATIC_REG1_ADDR};
        bins CH4_STATIC_REG2 = {`CH4_STATIC_REG2_ADDR};
        bins CH4_STATIC_REG3 = {`CH4_STATIC_REG3_ADDR};
        bins CH4_STATIC_REG4 = {`CH4_STATIC_REG4_ADDR};
        bins CH4_RESTRICT_REG = {`CH4_RESTRICT_REG_ADDR};
        bins CH4_READ_OFFSET_REG = {`CH4_READ_OFFSET_REG_ADDR};
        bins CH4_WRITE_OFFSET_REG = {`CH4_WRITE_OFFSET_REG_ADDR};
        bins CH4_FIFO_FULLNESS_REG = {`CH4_FIFO_FULLNESS_REG_ADDR};
        bins CH4_CMD_OUTS_REG = {`CH4_CMD_OUTS_REG_ADDR};
        bins CH4_CH_ENABLE_REG = {`CH4_CH_ENABLE_REG_ADDR};
        bins CH4_CH_START_REG = {`CH4_CH_START_REG_ADDR};
        bins CH4_CH_ACTIVE_REG = {`CH4_CH_ACTIVE_REG_ADDR};
        bins CH4_COUNT_REG = {`CH4_COUNT_REG_ADDR};
        bins CH4_INT_RAWSTAT_REG = {`CH4_INT_RAWSTAT_REG_ADDR};
        bins CH4_INT_CLEAR_REG = {`CH4_INT_CLEAR_REG_ADDR};
        bins CH4_INT_ENABLE_REG = {`CH4_INT_ENABLE_REG_ADDR};
        bins CH4_INT_STATUS_REG = {`CH4_INT_STATUS_REG_ADDR};
        bins CH5_CMD_REG0 = {`CH5_CMD_REG0_ADDR};
        bins CH5_CMD_REG1 = {`CH5_CMD_REG1_ADDR};
        bins CH5_CMD_REG2 = {`CH5_CMD_REG2_ADDR};
        bins CH5_CMD_REG3 = {`CH5_CMD_REG3_ADDR};
        bins CH5_STATIC_REG0 = {`CH5_STATIC_REG0_ADDR};
        bins CH5_STATIC_REG1 = {`CH5_STATIC_REG1_ADDR};
        bins CH5_STATIC_REG2 = {`CH5_STATIC_REG2_ADDR};
        bins CH5_STATIC_REG3 = {`CH5_STATIC_REG3_ADDR};
        bins CH5_STATIC_REG4 = {`CH5_STATIC_REG4_ADDR};
        bins CH5_RESTRICT_REG = {`CH5_RESTRICT_REG_ADDR};
        bins CH5_READ_OFFSET_REG = {`CH5_READ_OFFSET_REG_ADDR};
        bins CH5_WRITE_OFFSET_REG = {`CH5_WRITE_OFFSET_REG_ADDR};
        bins CH5_FIFO_FULLNESS_REG = {`CH5_FIFO_FULLNESS_REG_ADDR};
        bins CH5_CMD_OUTS_REG = {`CH5_CMD_OUTS_REG_ADDR};
        bins CH5_CH_ENABLE_REG = {`CH5_CH_ENABLE_REG_ADDR};
        bins CH5_CH_START_REG = {`CH5_CH_START_REG_ADDR};
        bins CH5_CH_ACTIVE_REG = {`CH5_CH_ACTIVE_REG_ADDR};
        bins CH5_COUNT_REG = {`CH5_COUNT_REG_ADDR};
        bins CH5_INT_RAWSTAT_REG = {`CH5_INT_RAWSTAT_REG_ADDR};
        bins CH5_INT_CLEAR_REG = {`CH5_INT_CLEAR_REG_ADDR};
        bins CH5_INT_ENABLE_REG = {`CH5_INT_ENABLE_REG_ADDR};
        bins CH5_INT_STATUS_REG = {`CH5_INT_STATUS_REG_ADDR};
        bins CH6_CMD_REG0 = {`CH6_CMD_REG0_ADDR};
        bins CH6_CMD_REG1 = {`CH6_CMD_REG1_ADDR};
        bins CH6_CMD_REG2 = {`CH6_CMD_REG2_ADDR};
        bins CH6_CMD_REG3 = {`CH6_CMD_REG3_ADDR};
        bins CH6_STATIC_REG0 = {`CH6_STATIC_REG0_ADDR};
        bins CH6_STATIC_REG1 = {`CH6_STATIC_REG1_ADDR};
        bins CH6_STATIC_REG2 = {`CH6_STATIC_REG2_ADDR};
        bins CH6_STATIC_REG3 = {`CH6_STATIC_REG3_ADDR};
        bins CH6_STATIC_REG4 = {`CH6_STATIC_REG4_ADDR};
        bins CH6_RESTRICT_REG = {`CH6_RESTRICT_REG_ADDR};
        bins CH6_READ_OFFSET_REG = {`CH6_READ_OFFSET_REG_ADDR};
        bins CH6_WRITE_OFFSET_REG = {`CH6_WRITE_OFFSET_REG_ADDR};
        bins CH6_FIFO_FULLNESS_REG = {`CH6_FIFO_FULLNESS_REG_ADDR};
        bins CH6_CMD_OUTS_REG = {`CH6_CMD_OUTS_REG_ADDR};
        bins CH6_CH_ENABLE_REG = {`CH6_CH_ENABLE_REG_ADDR};
        bins CH6_CH_START_REG = {`CH6_CH_START_REG_ADDR};
        bins CH6_CH_ACTIVE_REG = {`CH6_CH_ACTIVE_REG_ADDR};
        bins CH6_COUNT_REG = {`CH6_COUNT_REG_ADDR};
        bins CH6_INT_RAWSTAT_REG = {`CH6_INT_RAWSTAT_REG_ADDR};
        bins CH6_INT_CLEAR_REG = {`CH6_INT_CLEAR_REG_ADDR};
        bins CH6_INT_ENABLE_REG = {`CH6_INT_ENABLE_REG_ADDR};
        bins CH6_INT_STATUS_REG = {`CH6_INT_STATUS_REG_ADDR};
        bins CH7_CMD_REG0 = {`CH7_CMD_REG0_ADDR};
        bins CH7_CMD_REG1 = {`CH7_CMD_REG1_ADDR};
        bins CH7_CMD_REG2 = {`CH7_CMD_REG2_ADDR};
        bins CH7_CMD_REG3 = {`CH7_CMD_REG3_ADDR};
        bins CH7_STATIC_REG0 = {`CH7_STATIC_REG0_ADDR};
        bins CH7_STATIC_REG1 = {`CH7_STATIC_REG1_ADDR};
        bins CH7_STATIC_REG2 = {`CH7_STATIC_REG2_ADDR};
        bins CH7_STATIC_REG3 = {`CH7_STATIC_REG3_ADDR};
        bins CH7_STATIC_REG4 = {`CH7_STATIC_REG4_ADDR};
        bins CH7_RESTRICT_REG = {`CH7_RESTRICT_REG_ADDR};
        bins CH7_READ_OFFSET_REG = {`CH7_READ_OFFSET_REG_ADDR};
        bins CH7_WRITE_OFFSET_REG = {`CH7_WRITE_OFFSET_REG_ADDR};
        bins CH7_FIFO_FULLNESS_REG = {`CH7_FIFO_FULLNESS_REG_ADDR};
        bins CH7_CMD_OUTS_REG = {`CH7_CMD_OUTS_REG_ADDR};
        bins CH7_CH_ENABLE_REG = {`CH7_CH_ENABLE_REG_ADDR};
        bins CH7_CH_START_REG = {`CH7_CH_START_REG_ADDR};
        bins CH7_CH_ACTIVE_REG = {`CH7_CH_ACTIVE_REG_ADDR};
        bins CH7_COUNT_REG = {`CH7_COUNT_REG_ADDR};
        bins CH7_INT_RAWSTAT_REG = {`CH7_INT_RAWSTAT_REG_ADDR};
        bins CH7_INT_CLEAR_REG = {`CH7_INT_CLEAR_REG_ADDR};
        bins CH7_INT_ENABLE_REG = {`CH7_INT_ENABLE_REG_ADDR};
        bins CH7_INT_STATUS_REG = {`CH7_INT_STATUS_REG_ADDR};
        bins INT0_STATUS = {`INT0_STATUS_ADDR};
        bins CORE0_JOINT_MODE = {`CORE0_JOINT_MODE_ADDR};
        bins CORE0_PRIORITY = {`CORE0_PRIORITY_ADDR};
        bins CORE0_CH_START = {`CORE0_CH_START_ADDR};
        bins PERIPH_RX_CTRL = {`PERIPH_RX_CTRL_ADDR};
        bins PERIPH_TX_CTRL = {`PERIPH_TX_CTRL_ADDR};
        bins IDLE = {`IDLE_ADDR};
        bins USER_DEF_STATUS = {`USER_DEF_STATUS_ADDR};
        bins USER_CORE0_DEF_STATUS0 = {`USER_CORE0_DEF_STATUS0_ADDR};
        bins USER_CORE0_DEF_STATUS1 = {`USER_CORE0_DEF_STATUS1_ADDR};
	}
	WR_RD_CP: coverpoint tx.wr_rd;
	CROSS_ADDR_WR_RD: cross ADDR_CP,WR_RD_CP;
endgroup

function new(string name="",uvm_component parent);
	super.new(name,parent);
	apb_cg=new();
endfunction

function void build_phase(uvm_phase phase);
	super.build_phase(phase);
endfunction

function void write(apb_tx t);
	$cast(tx,t);
	apb_cg.sample();
endfunction
endclass
