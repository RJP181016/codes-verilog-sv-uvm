program test;
  
  `include "uvm_macros.svh"
  import uvm_pkg::*;
  `include "test.sv"
  
  initial run_test("new_test");
  
endprogram
