class eth_common;
endclass
