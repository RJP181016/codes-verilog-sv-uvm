`include "axi_intf.sv"
`include "axi_tx.sv"
`include "axi_slave.sv"
`include "axi_assertion.sv"
`include "axi_bfm.sv"
`include "axi_gen.sv"
`include "axi_mon.sv"
`include "axi_cov.sv"
`include "axi_env.sv"
`include "axi_tb.sv"
